
 module duck_game_logic

    (
        input  wire  clk,  // posedge active clock
        input  wire  rst,  // high-level active synchronous reset
        
        input  wire  [11:0] mouse_xpos, 
        input  wire  [11:0] mouse_ypos,
        input  wire  left_mouse,
        input  wire  right_mouse,
        input  wire  game_enable,

        input  wire  [11:0] duck_xpos,
        input  wire  [11:0] duck_ypos,

        output logic [2:0] bullets_in_magazine,
        output logic [5:0] bullets_left,
        output logic [6:0] my_score,
        output logic hunt_start,
        output logic show_reload_char
    );
    
    //------------------------------------------------------------------------------
    // local parameters
    //------------------------------------------------------------------------------
    localparam DUCK_HEIGHT = 60;
    localparam DUCK_WIDTH = 96;
    localparam STATE_BITS = 3; // number of bits used for state register

    // localparam COUNTDOWN    = 4000 * 65_000; // countdown value at start of the game T - 4000ms
    // localparam DEATH_TIME   = 2000 * 65_000; // time for duck fall after death T - 2000ms
    // localparam RELOAD_TIME  = 100 * 65_000; // time for reloading T - 100ms
    //FOR TESTS
    localparam COUNTDOWN    = 40; 
    localparam DEATH_TIME   = 20; 
    localparam RELOAD_TIME  = 1; 
    //------------------------------------------------------------------------------
    // local variables
    //------------------------------------------------------------------------------
    logic [2:0] bullets_in_magazine_nxt;
    logic [5:0] bullets_left_nxt;
    logic left_mouse_prev, left_mouse_posedge, right_mouse_posedge, right_mouse_prev;
    logic [31:0] delay_ms, delay_ms_nxt;
    logic [6:0] my_score_nxt;
    logic hunt_start_nxt, show_reload_char_nxt;
    
    enum logic [STATE_BITS-1 :0] {
        WAIT_FOR_START = 3'b000,
        HUNTING        = 3'b001,
        RELOADING      = 3'b010,
        DELAY          = 3'b011
    } state, state_nxt;
    
    //------------------------------------------------------------------------------
    // state sequential with synchronous reset
    //------------------------------------------------------------------------------
    always_ff @(posedge clk) begin : state_seq_blk
        if(rst)begin : state_seq_rst_blk
            state <= WAIT_FOR_START;
        end
        else begin : state_seq_run_blk
            state <= state_nxt;
        end
    end
    //------------------------------------------------------------------------------
    // next state logic
    //------------------------------------------------------------------------------
    always_comb begin : state_comb_blk
        case(state)
            WAIT_FOR_START: state_nxt = (game_enable) ? DELAY : WAIT_FOR_START;
            DELAY:          state_nxt = (delay_ms == 0) ? HUNTING : DELAY;
            HUNTING:
                if (right_mouse_posedge) 
                    state_nxt = RELOADING;
                else if (delay_ms == DEATH_TIME) 
                    state_nxt = DELAY;
                else 
                    state_nxt = HUNTING;

            RELOADING:      state_nxt = DELAY;
        endcase
    end
    //------------------------------------------------------------------------------
    // output register
    //------------------------------------------------------------------------------
    always_ff @(posedge clk) begin : out_reg_blk
        if(rst) begin : out_reg_rst_blk
            {bullets_in_magazine, bullets_left} <= 0;
            delay_ms <= COUNTDOWN;
            left_mouse_prev <= 0;
            right_mouse_prev <= 0;
            my_score <= 0;
            hunt_start <= 0;
            show_reload_char <= 0;
        end
        else begin : out_reg_run_blk
            bullets_in_magazine <= bullets_in_magazine_nxt;
            bullets_left <= bullets_left_nxt;
            delay_ms <= delay_ms_nxt;
            left_mouse_prev <= left_mouse;
            right_mouse_prev <= right_mouse;
            my_score <= my_score_nxt;
            hunt_start <= hunt_start_nxt;
            show_reload_char <= show_reload_char_nxt;
        end
    end
    //------------------------------------------------------------------------------
    // output logic
    //------------------------------------------------------------------------------
    always_comb begin : out_comb_blk
        left_mouse_posedge = (left_mouse == 1 && left_mouse_prev == 0);
        right_mouse_posedge = (right_mouse == 1 && right_mouse_prev == 0);
        case(state_nxt)
            WAIT_FOR_START: begin
                hunt_start_nxt = 0;
                delay_ms_nxt = COUNTDOWN;
                bullets_in_magazine_nxt = 3;
                bullets_left_nxt = 30;
                show_reload_char_nxt = 0;
                my_score_nxt = 0;
            end
            DELAY: begin
                hunt_start_nxt = 0;
                delay_ms_nxt = delay_ms - 1;
                bullets_in_magazine_nxt = bullets_in_magazine;
                bullets_left_nxt = bullets_left;
                show_reload_char_nxt = 0;
                my_score_nxt = my_score;
            end
            HUNTING: begin
                hunt_start_nxt = 1;
                delay_ms_nxt = delay_ms;
                bullets_in_magazine_nxt = bullets_in_magazine;
                bullets_left_nxt = bullets_left;
                show_reload_char_nxt = show_reload_char;
                my_score_nxt = my_score;

                if (left_mouse_posedge) begin
                    if (bullets_in_magazine > 0) begin
                        bullets_in_magazine_nxt = bullets_in_magazine - 1;
                        bullets_left_nxt = bullets_left - 1;
                        if (mouse_xpos >= duck_xpos && mouse_xpos <= duck_xpos + DUCK_WIDTH &&
                            mouse_ypos >= duck_ypos && mouse_ypos <= duck_ypos + DUCK_HEIGHT) begin
                            my_score_nxt = my_score + 1;
                            delay_ms_nxt = DEATH_TIME;
                        end
                    end else begin
                        show_reload_char_nxt = 1;
                    end
                end
            end

            RELOADING: begin
                hunt_start_nxt = 1;
                delay_ms_nxt = RELOAD_TIME;
                bullets_in_magazine_nxt = 3;
                bullets_left_nxt = bullets_left + bullets_in_magazine - 3;
                show_reload_char_nxt = 0;
                my_score_nxt = my_score;
            end
        endcase
    end
    
    endmodule
    