/**
 * San Jose State University
 * EE178 Lab #4
 * Author: prof. Eric Crabilla
 *
 * Modified by:
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Piotr Kaczmarczyk,
 * Łukasz Gąsecki
 * Oliwia Szewczyk
 * Description:
 * The project top module.
 */

module top_vga (
        input  logic clk65,
        input  logic rst,

        output logic vs,
        output logic hs,
        output logic [3:0] r,
        output logic [3:0] g,
        output logic [3:0] b,
        inout ps2_clk,
        inout ps2_data

    );

    timeunit 1ns;
    timeprecision 1ps;

     /**
     * Interface declarations
      */


    timing_if timing_if();
    vga_if background_if();
    vga_if draw_mouse_if();
    vga_if mouse_shape_if();
    vga_if game_if();


    /**
     * Local variables and signals
     */

    import vga_pkg::*;

    logic [11:0]xpos;
    logic [11:0]ypos;
    logic left_mouse, right_mouse;

    
    /**
     * Signals assignments
     */
    
    assign vs = game_if.vsync;
    assign hs = game_if.hsync;
    assign {r,g,b} = game_if.rgb;
    
    
    /**
     * Submodules instances
     */
    
    MouseCtl u_MouseCtl (
        .ps2_clk (ps2_clk),
        .ps2_data (ps2_data),
        .xpos (xpos),
        .ypos (ypos),
        .clk (clk65),
        .rst (rst),
        .value(12'b0),
        .setx('b0),
        .sety('b0),
        .setmax_x('b0),
        .setmax_y('b0),
        .new_event(),
        .zpos(),
        .left(left_mouse),
        .middle(),
        .right(right_mouse)
    );

    vga_timing u_vga_timing (
        .clk(clk65),
        .rst,

        .out(timing_if)
    );

    Game_Background u_game_background (
        .clk(clk65),
        .rst(rst),

        .in(timing_if),
        .out(background_if)
    );

    draw_mouse u_draw_mouse(
        .rst,   
        .clk(clk65),
        .xpos(xpos),
        .ypos(ypos),
        
        .in(mouse_shape_if),
        .out(draw_mouse_if)        
    );

    mouse_shape u_mouse_shape (
        .clk(clk65),
        .rst,
        .xpos (xpos),
        .ypos (ypos),
        .in(background_if),
        .out(mouse_shape_if)

    );

    top_game u_top_game (
        .clk(clk65),
        .rst(rst),
        .mouse_xpos(xpos),
        .mouse_ypos(ypos),
        .left_mouse(left_mouse),
        .right_mouse(right_mouse),

        .in(mouse_shape_if),
        .out(game_if)
    );

 
endmodule
